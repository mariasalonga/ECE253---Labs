module part1 (
    input logic Clock,
    input logic Enable,
    input logic Reset,
    output logic [7:0] CounterValue
);

module T_flip_flop (
                    input logic Clock,
                    

)